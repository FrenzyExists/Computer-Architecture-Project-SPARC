`timescale 1ns / 1ns

module alu_tester;

reg a;
reg b;

wire y;

mini_alu(
    
);

endmodule