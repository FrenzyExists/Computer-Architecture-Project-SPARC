


module sparc_fantastica(


);

endmodule