module condition_handler(
    input psr,
    input cwp, // Current Window Pointer
    output choose_branch
);

always@(*) begin
    if()
    
    endif
end

endmodule